module randomm(clk, choose, en, data_in, Q, seg0, seg1);
	input [2:0] choose;
	input en;
	input [7:0] data_in;
	input clk;
	output reg [7:0] Q;
	reg inone;
	output reg [6:0] seg0;
	output reg [6:0] seg1;
	reg [3:0] Qh;
	reg [3:0] Ql;
	reg replace = 0;
	reg out1;
	reg out2;
	always @(posedge clk)
	begin
		if(en)
			begin
				case(choose)
				0:Q = 0;
				1:Q = data_in;
				2:Q = {replace, Q[7:1]};
				3:Q = {Q[6:0], replace};
				4:Q = {Q[7], Q[7:1]};
				5:begin out1 = Q[4] ^ Q[3] ^ Q[2] ^ Q[0]; out2 = ~(Q[7] | Q[6] | Q[5] | Q[4] | Q[3] | Q[2] | Q[1]); inone = out1 ^ out2; Q = {inone, Q[7:1]}; end
				6:Q = {Q[0], Q[7:1]};
				7:Q = {Q[6:0], Q[7]};
				endcase
			end
		else
		begin
			Q = 0;
		end
		Qh = Q[7:4];
		Ql = Q[3:0];
		case(Qh)
		0: seg1 = 7'b1000000;
		1: seg1 = 7'b1111001;
		2: seg1 = 7'b0100100;
		3: seg1 = 7'b0110000;
		4: seg1 = 7'b0011001;
		5: seg1 = 7'b0010010;
		6: seg1 = 7'b0000010;
		7: seg1 = 7'b1111000;
		8: seg1 = 7'b0000000;
		9: seg1 = 7'b0010000;
		10: seg1 = 7'b0001000;
		11: seg1 = 7'b0000011;
		12: seg1 = 7'b1000110;
		13: seg1 = 7'b0100001;
		14: seg1 = 7'b0000110;
		15: seg1 = 7'b0001110;
		endcase

		case(Ql)
		0: seg0 = 7'b1000000;
		1: seg0 = 7'b1111001;
		2: seg0 = 7'b0100100;
		3: seg0 = 7'b0110000;
		4: seg0 = 7'b0011001;
		5: seg0 = 7'b0010010;
		6: seg0 = 7'b0000010;
		7: seg0 = 7'b1111000;
		8: seg0 = 7'b0000000;
		9: seg0 = 7'b0010000;
		10: seg0 = 7'b0001000;
		11: seg0 = 7'b0000011;
		12: seg0 = 7'b1000110;
		13: seg0 = 7'b0100001;
		14: seg0 = 7'b0000110;
		15: seg0 = 7'b0001110;
		endcase
	end
endmodule